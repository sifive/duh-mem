module ram1 (

);

endmodule
